/****************************************************************************
 * Copyright (c) 2009 by Focus Robotics. All rights reserved.
 *
 * This program is an unpublished work fully protected by the United States 
 * copyright laws and is considered a trade secret belonging to the copyright
 * holder. No part of this design may be reproduced stored in a retrieval 
 * system, or transmitted, in any form or by any means, electronic, 
 * mechanical, photocopying, recording, or otherwise, without prior written 
 * permission of Focus Robotics, Inc.
 *
 * Proprietary and Confidential
 *
 * Created By   :  Andrew Worcester
 * Creation_Date:  Tue Mar 10 2009
 * 
 * Brief Description:
 * 
 * Functionality:
 * 
 * Issues:
 * 
 * Limitations:
 * 
 * Testing:
 * 
 * Synthesis:
 * 
 ******************************************************************************/

module fric_switch_8port
  (
   clk,
   rst,
   fric_in0,
   fric_out0,
   fric_in1,
   fric_out1,
   fric_in2,
   fric_out2,
   fric_in3,
   fric_out3,
   fric_in4,
   fric_out4,
   fric_in5,
   fric_out5,
   fric_in6,
   fric_out6,
   fric_in7,
   fric_out7
   );

   // In/Out declarations
   input           clk;
   input 	   rst;
   input [7:0] 	   fric_in0;
   output [7:0]    fric_out0;
   input [7:0] 	   fric_in1;
   output [7:0]    fric_out1;
   input [7:0] 	   fric_in2;
   output [7:0]    fric_out2;
   input [7:0] 	   fric_in3;
   output [7:0]    fric_out3;
   input [7:0] 	   fric_in4;
   output [7:0]    fric_out4;
   input [7:0] 	   fric_in5;
   output [7:0]    fric_out5;
   input [7:0] 	   fric_in6;
   output [7:0]    fric_out6;
   input [7:0] 	   fric_in7;
   output [7:0]    fric_out7;

   // Parameters

   // Regs and Wires

   // RTL or Instances

   /****************************************************************************
    * Subblock
    * 
    * Inputs:
    * 
    * Outputs:
    * 
    * Todo/Fixme:
    * 
    */
   

endmodule // fric_switch_8port





